package rv;
  typedef enum logic [10:0] {
    LUI   = 11'bx_xxx_0110111,
    AUIPC = 11'bx_xxx_0010111,
    JAL   = 11'bx_xxx_1101111,
    JALR  = 11'bx_000_1100111,
    BEQ   = 11'bx_000_1100011,
    BNE   = 11'bx_001_1100011,
    BLT   = 11'bx_100_1100011,
    BGE   = 11'bx_101_1100011,
    BLTU  = 11'bx_110_1100011,
    BGEU  = 11'bx_111_1100011,
    LB    = 11'bx_000_0000011,
    LH    = 11'bx_001_0000011,
    LW    = 11'bx_010_0000011,
    LBU   = 11'bx_100_0000011,
    LHU   = 11'bx_101_0000011,
    SB    = 11'bx_000_0100011,
    SH    = 11'bx_001_0100011,
    SW    = 11'bx_010_0100011,
    ADDI  = 11'bx_000_0010011,
    SLTI  = 11'bx_000_0010011,
    SLTIU = 11'bx_011_0010011,
    XORI  = 11'bx_100_0010011,
    ORI   = 11'bx_110_0010011,
    ANDI  = 11'bx_111_0010011,
    SLLI  = 11'b0_001_0010011,
    SRLI  = 11'b0_101_0010011,
    SRAI  = 11'b1_101_0010011,
    ADD   = 11'b0_000_0110110,
    SUB   = 11'b1_000_0110110,
    SLL   = 11'b0_001_0110011,
    SLT   = 11'b0_010_0110011,
    SLTU  = 11'b0_011_0110011,
    XOR   = 11'b0_100_0110011,
    SRL   = 11'b0_101_0110011,
    SRA   = 11'b1_101_0110011,
    OR    = 11'b0_110_0110011,
    AND   = 11'b0_111_0110011
  } RV32_INSTRUCTION;
endpackage
